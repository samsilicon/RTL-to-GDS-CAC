/home/sameer25145/Desktop/CAC_Project_Part2/IN/lef/gsclib090_translated_ref.lef